library verilog;
use verilog.vl_types.all;
entity full_adder_tb is
end full_adder_tb;
